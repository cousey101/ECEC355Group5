LIBRARY ieee;
USE ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use ieee.numeric_std.all;

entity 1bALU is
port(
	a,b,aInv,bInv,oper,less,cIn:in std_logic_vector(1 downto 0);
	result,cOut:out std_logic_vector(1 downto 0));
  
end 1bALU;

ARCHITECTURE beh of 1bALU is
begin
end beh;